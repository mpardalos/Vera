module add(input reg [31:0] x, input reg [31:0] y, output wire [31:0] out);
   assign out = x + y;
endmodule // add
