module Mult(input in1, input in2, output out);
   wire [31:0] in1;
   wire [31:0] in2;
   wire [31:0] out;

   assign out = in1 + (0 + in2);
endmodule // Shift
