module add(output reg [31:0] out);
   assign out = 1 + 2;
endmodule // add
